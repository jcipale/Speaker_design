subwoofer-zobel
*----------------------------------------------
*	GNUCAP - NETLIST
.options OUT=120 
*------------- Models -------------------------
*------------- Circuit Description-------------
R_Rz1 4 0 6.2
R_Spk1 6 0 
V_V1 3 0 dc 0.0 ac 1.0 sin(0.0 1.0 1.0 0 0)
R_R1 5 6 6.2
L_L2 1 5 1H
C_C1 2 1 1u IC=0
C_Cz1 1 4 0.0156u IC=0
L_L1 3 2 15.9m

*----------------------------------------------
* Analysis Requests
*----------------------------------------------
*.print tran  v(6)
.tran 0 0.005 5e-05
.print op v(nodes)
.op
.end
